module andGate(in0,in1,in2,out);
input in0,in1,in2;
output out;

assign out = in0&in1&in2;
endmodule